
module data_mem(input [31:0] addr, input [31:0] writeData, input memRead, input memWrite, output reg [31:0]readData);
	
	reg [32:0] ram [15:0];
	initial 
	begin 
			ram[0] = 32'b00000000000000000000000000000000;  
            ram[1] = 32'b00000000000000000000000000000001; 
            ram[2] = 32'b00000000000000000000000000000010;  
            ram[3] = 32'b00000000000000000000000000000011;  
            ram[4] = 32'b00000000000000000000000000000100;  
            ram[5] = 32'b00000000000000000000000000000101;
            ram[6] = 32'b00000000000000000000000000000111;  
            ram[7] = 32'b00000000000000000000000000001000; 
            ram[8] = 32'b00000000000000000000000000000000;  
            ram[9] = 32'b00000000000000000000000000000000; 
            ram[10] = 32'b00000000000000000000000000000000;  
            ram[11] = 32'b00000000000000000000000000000000;  
            ram[12] = 32'b00000000000000000000000000000000;
            ram[13] = 32'b00000000000000000000000000000000;  
            ram[14] = 32'b00000000000000000000000000000000;  
            ram[15] = 32'b00000000000000000000000000000000;
	end 
	always@ (addr,writeData,memRead,memWrite) begin
	
	 readData =  memRead ? ram[addr] : 32'b0 ;

	if (memWrite)
 		ram[addr] <= writeData;
	end
endmodule