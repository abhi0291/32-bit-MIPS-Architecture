
module instr_mem(input [31:0] addr, output [31:0] instr); 
	reg [32:0] rom[15:0];
	assign instr =  addr < 16 ? rom[addr[31:0]] : 32'b0 ;
	initial 
		begin 
		
		/*rom[0] = 32'b00000001010010110100100000100010;  //sub t1 t2 t3;
                rom[1] = 32'b00010010101101100000000000000010; 	//beq s5 s6 0x2;
                rom[2] = 32'b00000001100011010101100000100000;  //add t3 t4 t5;
                rom[3] = 32'b00000001101011100110000000100000;  //add t4 t5 t6;
                rom[4] = 32'b00000001110011110110100000100000;  //add t5 t6 t7;
                rom[5] = 32'b10001110010100010000000000000010;	//lw s1 0x2 s2;
                rom[6] = 32'b00000000000000000000000000000000;  
                rom[7] = 32'b00000000000000000000000000000000;  
                rom[8] = 32'b00000000000000000000000000000000;  
                rom[9] = 32'b00000000000000000000000000000000; 
                rom[10] = 32'b00000000000000000000000000000000;  
                rom[11] = 32'b00000000000000000000000000000000;  
                rom[12] = 32'b00000000000000000000000000000000;
                rom[13] = 32'b00000000000000000000000000000000;  
                rom[14] = 32'b00000000000000000000000000000000;
				rom[15] = 32'b00000000000000000000000000000000;*/
				rom[0] = 32'b10001110010100010000000000000010;  //sub t1 t2 t3;
                rom[1] = 32'b00000000000000000000000000000000; 	//beq s5 s6 0x2;
                rom[2] = 32'b00000000000000000000000000000000;  //add t3 t4 t5;
                rom[3] = 32'b00000000000000000000000000000000;  //add t4 t5 t6;
                rom[4] = 32'b00000000000000000000000000000000;  //add t5 t6 t7;
                rom[5] = 32'b100000000000000000000000000000000;	//lw s1 0x2 s2;
                rom[6] = 32'b00000000000000000000000000000000;  
                rom[7] = 32'b00000000000000000000000000000000;  
                rom[8] = 32'b00000000000000000000000000000000;  
                rom[9] = 32'b00000000000000000000000000000000; 
                rom[10] = 32'b00000000000000000000000000000000;  
                rom[11] = 32'b00000000000000000000000000000000;  
                rom[12] = 32'b00000000000000000000000000000000;
                rom[13] = 32'b00000000000000000000000000000000;  
                rom[14] = 32'b00000000000000000000000000000000;
				rom[15] = 32'b00000000000000000000000000000000;
		
		end 
	
endmodule