module registers_file ( input reg_write , input [4:0]  read_reg1 , input [4:0] read_reg2, input [4:0] write_reg , input [31:0] write_data
			, output reg [31:0] read_data1 , output reg [31:0] read_data2 );
	
	reg [31:0] registors[31:0];
	
	initial begin 

	registors[0] <= 32'b00000000000000000000000000000000; //$0
	registors[1] <= 32'b00000000000000000000000000000000;
	registors[2] <= 32'b00000000000000000000000000000000;
	registors[3] <= 32'b00000000000000000000000000000000;
	registors[4] <= 32'b00000000000000000000000000000000;
	registors[5] <= 32'b00000000000000000000000000000000;
	registors[6] <= 32'b00000000000000000000000000000000;
	registors[7] <= 32'b00000000000000000000000000000000;
	registors[8] <= 32'b00000000000000000000000000000000; //$t0
	registors[9] <= 32'b00000000000000000000000000000001;
	registors[10] <= 32'b00000000000000000000000000000010;
	registors[11] <= 32'b00000000000000000000000000000011;
	registors[12] <= 32'b00000000000000000000000000000100;
	registors[13] <= 32'b00000000000000000000000000000101;
	registors[14] <= 32'b00000000000000000000000000000110;
	registors[15] <= 32'b00000000000000000000000000000111; //$t7
	registors[16] <= 32'b00000000000000000000000000001000; //$s0
	registors[17] <= 32'b00000000000000000000000000001001;
	registors[18] <= 32'b00000000000000000000000000000001;
	registors[19] <= 32'b00000000000000000000000000001011;
	registors[20] <= 32'b00000000000000000000000000001100;
	registors[21] <= 32'b00000000000000000000000000001101;
	registors[22] <= 32'b00000000000000000000000000001101;
	registors[23] <= 32'b00000000000000000000000000001111; //$s7
	registors[24] <= 32'b00000000000000000000000000000000;
	registors[25] <= 32'b00000000000000000000000000000000;
	registors[26] <= 32'b00000000000000000000000000000000;
	registors[27] <= 32'b00000000000000000000000000000000;
	registors[28] <= 32'b00000000000000000000000000000000;
	registors[29] <= 32'b00000000000000000000000000000000;
	registors[30] <= 32'b00000000000000000000000000000000;
	registors[31] <= 32'b00000000000000000000000000000000;

	end 	

	always @( reg_write , read_reg1 , read_reg2 , write_reg , write_data ) begin
	if (reg_write) begin
		registors[write_reg] <= write_data;
		end
	read_data1 <= registors[read_reg1];
	read_data2 <= registors[read_reg2];
	end
			 
endmodule